module ulaaux (
    input wire [31:0] A,
    input wire [31:0] B,
    input wire [1:0] ulaaux_control, // Operações a ser definidas
    output wire ulaux_out,
    output wire SPECIAL
);


endmodule